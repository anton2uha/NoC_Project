
//virtual channel allocator
module VCA (
	input wire [63:0] creditsIn, in_northBuf, in_eastBuf, in_southBuf, in_westBuf,
	output wire [63:0] creditsOut, out_northBuf, out_eastBuf, out_southBuf, out_westBuf
	
);




endmodule