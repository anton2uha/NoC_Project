
module Buffer (
	input wire [63:0] dataIn, in_VCA, in_RC, in_CBA,
	output wire [63:0]out_CBS, out_VCA, out_RC, out_CBA

);






endmodule
