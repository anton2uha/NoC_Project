
module CrossBarSwitch (
	input wire [63:0] northBuf, eastBuf, southBuf, westBuf, in_CBA,
	
	output wire [63:0] northOut, eastOut, southOut, westOut, out_CBA

);



endmodule