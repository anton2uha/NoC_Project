
// route computation unit
module RC (
	input wire [63:0] in_northBuf, in_eastBuf, in_southBuf, in_westBuf,
	output wire [63:0] out_northBuf, out_eastBuf, out_southBuf, out_westBuf
);



endmodule