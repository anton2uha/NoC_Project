
//processing unit
module PE (
	input wire [63:0] routerIn,
	output wire [63:0] routerOut
);




endmodule